//======================================================================
//
// sha256_w_mem_regs.v
// -------------------
// The W memory. This includes functionality to expand the block
// into 64 words. This is the old version based on separate registers.
// This version is saved as a loose module to be used if the
// synthesis tool is unable to do proper mapping of the array
// based implementation.
//
//
// Copyright (c) 2013 Secworks Sweden AB
// All rights reserved.
// 
// Redistribution and use in source and binary forms, with or 
// without modification, are permitted provided that the following 
// conditions are met: 
// 
// 1. Redistributions of source code must retain the above copyright 
//    notice, this list of conditions and the following disclaimer. 
// 
// 2. Redistributions in binary form must reproduce the above copyright 
//    notice, this list of conditions and the following disclaimer in 
//    the documentation and/or other materials provided with the 
//    distribution. 
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS 
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT 
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS 
// FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE 
// COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, 
// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, 
// BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER 
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, 
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) 
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF 
// ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//======================================================================

module sha256_w_mem(
                    input wire           clk,
                    input wire           reset_n,

                    input wire [511 : 0] block,

                    input wire           init,
                    input wire           next,
                    output wire [31 : 0] w
                   );

  
  //----------------------------------------------------------------
  // Internal constant and parameter definitions.
  //----------------------------------------------------------------
  parameter CTRL_IDLE   = 0;
  parameter CTRL_UPDATE = 1;
  
  
  //----------------------------------------------------------------
  // Registers including update variables and write enable.
  //----------------------------------------------------------------
  reg [31 : 0] w_mem [0 : 15];
  
  reg [5 : 0] w_ctr_reg;
  reg [5 : 0] w_ctr_new;
  reg         w_ctr_we;
  reg         w_ctr_inc;
  reg         w_ctr_rst;
  
  reg [1 : 0]  sha256_w_mem_ctrl_reg;
  reg [1 : 0]  sha256_w_mem_ctrl_new;
  reg          sha256_w_mem_ctrl_we;
  
  
  //----------------------------------------------------------------
  // Wires.
  //----------------------------------------------------------------
  reg [31 : 0] w_tmp;
  reg [31 : 0] w_new;
  
  reg w_update;
  reg mem_update;
  
  
  //----------------------------------------------------------------
  // Concurrent connectivity for ports etc.
  //----------------------------------------------------------------
  assign w = w_tmp;
  
  
  //----------------------------------------------------------------
  // reg_update
  // Update functionality for all registers in the core.
  // All registers are positive edge triggered with synchronous
  // active low reset. All registers have write enable.
  //----------------------------------------------------------------
  always @ (posedge clk)
    begin : reg_update
      if (!reset_n)
        begin
          w_ctr_reg             <= 6'h00;
          sha256_w_mem_ctrl_reg <= CTRL_IDLE;
        end
      else
        begin
          if (init)
            begin
              w_mem[00] <= block[511 : 480];
              w_mem[01] <= block[479 : 448];
              w_mem[02] <= block[447 : 416];
              w_mem[03] <= block[415 : 384];
              w_mem[04] <= block[383 : 352];
              w_mem[05] <= block[351 : 320];
              w_mem[06] <= block[319 : 288];
              w_mem[07] <= block[287 : 256];
              w_mem[08] <= block[255 : 224];
              w_mem[09] <= block[223 : 192];
              w_mem[10] <= block[191 : 160];
              w_mem[11] <= block[159 : 128];
              w_mem[12] <= block[127 :  96];
              w_mem[13] <= block[95  :  64];
              w_mem[14] <= block[63  :  32];
              w_mem[15] <= block[31  :   0];
            end
          else if (mem_update)
            begin
              w_mem[00] <= w_mem[01];
              w_mem[01] <= w_mem[02];
              w_mem[02] <= w_mem[03];
              w_mem[03] <= w_mem[04];
              w_mem[04] <= w_mem[05];
              w_mem[05] <= w_mem[06];
              w_mem[06] <= w_mem[07];
              w_mem[07] <= w_mem[08];
              w_mem[08] <= w_mem[09];
              w_mem[09] <= w_mem[10];
              w_mem[10] <= w_mem[11];
              w_mem[11] <= w_mem[12];
              w_mem[12] <= w_mem[13];
              w_mem[13] <= w_mem[14];
              w_mem[14] <= w_mem[15];
              w_mem[15] <= w_new;
            end
          
          if (w_ctr_we)
            begin
              w_ctr_reg <= w_ctr_new;
            end
          
          if (sha256_w_mem_ctrl_we)
            begin
              sha256_w_mem_ctrl_reg <= sha256_w_mem_ctrl_new;
            end
        end
    end // reg_update

  
  //----------------------------------------------------------------
  // external_addr_mux
  //
  // Mux for the external read operation. This is where we exract
  // the W variable.
  //----------------------------------------------------------------
  always @*
    begin : external_addr_mux
      if (w_ctr_reg < 16)
        begin
          w_tmp      = w_mem[w_ctr_reg[3 : 0]];
          mem_update = 0;
        end
      else
        begin
          w_tmp      = w_new;
          mem_update = 1;
        end
    end // external_addr_mux
  

  //----------------------------------------------------------------
  // w_new_logic
  //
  // Logic that calculates the next value to be inserted into
  // the sliding window of the memory.
  //----------------------------------------------------------------
  always @*
    begin : w_new_logic
      reg [31 : 0] w_0;
      reg [31 : 0] w_1;
      reg [31 : 0] w_9;
      reg [31 : 0] w_14;
      reg [31 : 0] d0;
      reg [31 : 0] d1;

      w_0  = w_mem[0];
      w_1  = w_mem[1];
      w_9  = w_mem[9];
      w_14 = w_mem[14];

      d0 = {w_1[6  : 0], w_1[31 :  7]} ^ 
           {w_1[17 : 0], w_1[31 : 18]} ^ 
           {3'b000, w_1[31 : 3]};
      
      d1 = {w_14[16 : 0], w_14[31 : 17]} ^ 
           {w_14[18 : 0], w_14[31 : 19]} ^ 
           {10'b0000000000, w_14[31 : 10]};
      
      w_new = d1 + w_9 + d0 + w_0;
    end // w_new_logic
  
  
  //----------------------------------------------------------------
  // w_ctr
  // W schedule adress counter. Counts from 0x10 to 0x3f and
  // is used to expand the block into words.
  //----------------------------------------------------------------
  always @*
    begin : w_ctr
      w_ctr_new = 0;
      w_ctr_we  = 0;
      
      if (w_ctr_rst)
        begin
          w_ctr_new = 6'h00;
          w_ctr_we  = 1;
        end

      if (w_ctr_inc)
        begin
          w_ctr_new = w_ctr_reg + 6'h01;
          w_ctr_we  = 1;
        end
    end // w_ctr

  
  //----------------------------------------------------------------
  // sha256_w_mem_fsm
  // Logic for the w shedule FSM.
  //----------------------------------------------------------------
  always @*
    begin : sha256_w_mem_fsm
      w_ctr_rst = 0;
      w_ctr_inc = 0;
      w_update  = 0;
      
      sha256_w_mem_ctrl_new = CTRL_IDLE;
      sha256_w_mem_ctrl_we  = 0;
      
      case (sha256_w_mem_ctrl_reg)
        CTRL_IDLE:
          begin
            if (init)
              begin
                w_ctr_rst             = 1;
                sha256_w_mem_ctrl_new = CTRL_UPDATE;
                sha256_w_mem_ctrl_we  = 1;
              end
          end
        
        CTRL_UPDATE:
          begin
            if (next)
              begin
                w_update  = 1;
                w_ctr_inc = 1;
              end
            
            if (w_ctr_reg == 6'h3f)
              begin
                sha256_w_mem_ctrl_new = CTRL_IDLE;
                sha256_w_mem_ctrl_we  = 1;
              end
          end
      endcase // case (sha256_ctrl_reg)
    end // sha256_ctrl_fsm

endmodule // sha256_w_mem

//======================================================================
// sha256_w_mem.v
//======================================================================
